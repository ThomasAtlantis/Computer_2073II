library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
entity rom is
	port(
		enrom, romin: in std_logic;
		rom_address: in std_logic_vector(7 downto 0);
		rom_data: out std_logic_vector(7 downto 0)
	);
end entity rom;
architecture behave of rom is
type t_rom is array(0 to 63) of std_logic_vector(7 downto 0);
constant inner_data: t_rom := (
"00001000", "00001111", "00001001", "00000011", "01101100", "00000001", "10010100", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --rom   8 to  15
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --rom  16 to  23
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --rom  24 to  31
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --32 to 39
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --40 to 47
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --48 to 55
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000"  --56 to 63
--"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --64 to 71
--"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --72 to 79
--"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --80 to 87
--"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --88 to 95
--"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --96 to 103
--"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --104 to 111
--"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --112 to 119
--"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --120 to 127
--"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --128 to 135
--"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --136 to 143
--"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --144 to 151
--"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --152 to 159
--"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --160 to 167
--"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --168 to 175
--"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --176 to 183
--"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --184 to 191
--"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --192 to 199
--"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --200 to 207
--"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --208 to 215
--"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --216 to 223
--"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --224 to 231
--"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --232 to 239
--"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --240 to 247
--"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000"  --248 to 255
);
signal rom_address_latch: std_logic_vector(7 downto 0) := (others => '0');
begin
	process(romin)
	begin
		if (romin'event and romin = '1') then
			rom_address_latch <= rom_address;
		else 
			rom_address_latch <= rom_address_latch;
		end if;
	end process;
	rom_data <= inner_data(CONV_INTEGER(rom_address_latch)) when enrom = '1' else (others => 'Z');
end behave;